library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_unsigned.ALL;
USE IEEE.numeric_std.ALL;

entity orb is

generic
(
    pairs_num : integer:=64;
    delay_clk:integer:=5

);


port(
    clk : in std_logic;
    rst : in std_logic;	
    kp_en : in std_logic;
    save_en : in std_logic;
    video_clk      : in std_logic;
    vga_hs_cnt : in integer range 0 to 857;
    vga_vs_cnt : in integer range 0 to 524;
--    pepiclk  : out integer;
    BOUT_1 : out std_logic_vector(83 downto 0);
    --pepi: OUT std_logic_vector(0 downto 0);
    ping_pong_out_2_out : out std_logic_vector(7 downto 0);
    video_data : in std_logic_vector(7 downto 0);
    TRACKORB : IN std_logic_vector(39 downto 0);
    TRACKX : IN integer;
    TRACKY : IN integer;
    TRACKSQ : IN integer
 );


end orb;
  
architecture Behavioral of orb is

    
    type   array_type is array (integer range -4 to 4,integer range -4 to 4) of std_logic_vector (7 downto 0); 
    signal centroid_array   : array_type ;
    signal centroid_array_1 : array_type ;
    signal centroid_array_2 : array_type ;
    signal centroid_array_3 : array_type ;
    -- signal centroid_reg     : array_type ;
    
    signal	centroid_x_out  : signed (14 downto 0); 	
    signal	centroid_y_out  : signed (14 downto 0); 	

    signal	centroid_angle  : integer range 0 to 360;
    signal	angle_range     : integer range 0 to 11;


    signal  brief_array : array_type;
    signal	x_out :  STD_LOGIC_VECTOR(17 downto 0);
    signal	y_out :  STD_LOGIC_VECTOR(17 downto 0);
    signal	z_out :  STD_LOGIC_VECTOR(7 downto 0);
    
    signal ping_pong_out_8, ping_pong_out_7, ping_pong_out_6, ping_pong_out_5 : std_logic_vector(7 downto 0);
    signal ping_pong_out_4, ping_pong_out_3, ping_pong_out_2 ,ping_pong_out_1 : std_logic_vector(7 downto 0);
    
    signal brief_code : std_logic_vector(63 downto 0);

    type   kn_delay is array(integer range 0 to (delay_clk-1))of std_logic;
    signal kn_stage : kn_delay;
    
    type   cnt_delay is array(integer range 0 to (delay_clk-1))of std_logic_vector(9 downto 0);
    signal h_cnt_delay, v_cnt_delay : cnt_delay ;

    signal save       : std_logic_vector(127 downto 0);

    signal dina_1     : std_logic_vector( 83 downto 0);
    signal addra_1    : std_logic_vector( 7 downto 0);
    signal wea_1      : std_logic_vector( 0 downto 0);

    signal dina_2     : std_logic_vector( 83 downto 0);
    signal addra_2    : std_logic_vector( 7 downto 0);
    signal wea_2      : std_logic_vector( 0 downto 0);

    signal save_cnt_1 : std_logic_vector( 7 downto 0);
    signal save_cnt_2 : std_logic_vector( 7 downto 0);

--    signal  h,v,X1,Y1,X2,Y2,TRACKX,TRACKY : integer;
    --------------------------------------------------------- table
    
    --128�I�� �d��
    type pairs_table is ARRAY(integer range  0 to  (pairs_num-1),integer range 0 to 12) of integer range -4 to  4;
    
    Constant y1_sin_pairs : pairs_table := 
    -- y1 sin
    --0     30     60     90    120    150    180    210    230    270    300    330    360
    --0      1      2      3      4      5      6      7      8      9     10     11     12
    (
    ( 0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0 ),
    ( 0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0 ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0 ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0 ),
    ( 0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0 ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0 ),
    ( 0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0 ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0 ),
    ( 0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0 ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0 ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0 ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0 ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0 ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0 ),
    ( 0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0 ),
    ( 0,     2,     3,     4,     3,     2,     0,    -2,    -3,    -4,    -3,    -2,     0 ),
    ( 0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0 ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0 ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0 ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0 ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0 ),
    ( 0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0 ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0 ),
    ( 0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0 ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0 ),
    ( 0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0 ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0 ),
    ( 0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0 ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0 ),
    ( 0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0 ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0 ),
    ( 0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0 ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0 ),
    ( 0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0 ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0 ),
    ( 0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0 ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0 ),
    ( 0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0 ),
    ( 0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0 ),
    ( 0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0 ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0 ),
    ( 0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0 ),
    ( 0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0 ),
    ( 0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0 ),
    ( 0,    -2,    -3,    -4,    -3,    -2,     0,     2,     3,     4,     3,     2,     0 ),
    ( 0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0 ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0 ),
    ( 0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0 ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0 ),
    ( 0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0 ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0 ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0 ),
    ( 0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0 )
    );

    Constant x1_sin_pairs : pairs_table := 
    -- x1 sin
    (
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0 ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0 ),
    ( 0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0 ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0 ),
    ( 0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0 ),
    ( 0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0 ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0 ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0 ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0 ),
    ( 0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0 ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0 ),
    ( 0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0 ),
    ( 0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0 ),
    ( 0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0 ),
    ( 0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0 ),
    ( 0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0 ),
    ( 0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0 ),
    ( 0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0 ),
    ( 0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0 ),
    ( 0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0 ),
    ( 0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0 ),
    ( 0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0 ),
    ( 0,     2,     3,     4,     3,     2,     0,    -2,    -3,    -4,    -3,    -2,     0 ),
    ( 0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0 ),
    ( 0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0 ),
    ( 0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0 ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0 ),
    ( 0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0 ),
    ( 0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0 ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0 ),
    ( 0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0 ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0 ),
    ( 0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0 ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0 ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0 ),
    ( 0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0 ),
    ( 0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0 ),
    ( 0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0 ),
    ( 0,    -2,    -3,    -4,    -3,    -2,     0,     2,     3,     4,     3,     2,     0 ),
    ( 0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0 ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0 ),
    ( 0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0 ),
    ( 0,     2,     3,     4,     3,     2,     0,    -2,    -3,    -4,    -3,    -2,     0 ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0 ),
    ( 0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0 ),
    ( 0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0 ),
    ( 0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0 ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0 ),
    ( 0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0 ),
    ( 0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0 ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0 ),
    ( 0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0 ),
    ( 0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0 ),
    ( 0,     2,     3,     4,     3,     2,     0,    -2,    -3,    -4,    -3,    -2,     0 ),
    ( 0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0 ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0 ),
    ( 0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0 ),
    ( 0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0 )
    );

    Constant y1_cos_pairs : pairs_table := 
    --y1 cos
    (
    ( 3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3  ),
    ( 3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3  ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( 3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3  ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3 ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1  ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( 1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1  ),
    ( 4,     3,     2,     0,    -2,    -3,    -4,    -3,    -2,     0,     2,     3,     4  ),
    ( -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2 ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3  ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2 ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( 3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3  ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3 ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2 ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3 ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2 ),
    ( 1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1  ),
    ( -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3 ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3 ),
    ( -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2 ),
    ( -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2 ),
    ( -4,    -3,    -2,     0,     2,     3,     4,     3,     2,     0,    -2,    -3,    -4 ),
    ( 3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3  ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3 ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3 ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2 )
    );
    
    Constant x1_cos_pairs : pairs_table := 
    --x1 cos
    (
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( 1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1  ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( 3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3  ),
    ( 3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3  ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2 ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( 3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3  ),
    ( 3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1  ),
    ( 1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1  ),
    ( 1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1  ),
    ( -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3 ),
    ( 1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1  ),
    ( -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2 ),
    ( -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3 ),
    ( -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3 ),
    ( -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2 ),
    ( 4,     3,     2,     0,    -2,    -3,    -4,    -3,    -2,     0,     2,     3,     4  ),
    ( -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2 ),
    ( -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1  ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3 ),
    ( 1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1  ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2 ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2 ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2 ),
    ( -4,    -3,    -2,     0,     2,     3,     4,     3,     2,     0,    -2,    -3,    -4 ),
    ( 3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3  ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( 1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1  ),
    ( 4,     3,     2,     0,    -2,    -3,    -4,    -3,    -2,     0,     2,     3,     4  ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( 1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1  ),
    ( -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2 ),
    ( -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2 ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( 1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1  ),
    ( -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2 ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2 ),
    ( 1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1  ),
    ( 4,     3,     2,     0,    -2,    -3,    -4,    -3,    -2,     0,     2,     3,     4  ),
    ( -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2 ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( 3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3  ),
    ( -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3 )
    );
    
    Constant y2_sin_pairs : pairs_table := 
    -- y2 sin
    (
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0  ),
    ( 0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0  ),
    ( 0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0  ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0  ),
    ( 0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0  ),
    ( 0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0  ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0  ),
    ( 0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0  ),
    ( 0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0  ),
    ( 0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0  ),
    ( 0,     2,     3,     4,     3,     2,     0,    -2,    -3,    -4,    -3,    -2,     0  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0  ),
    ( 0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0  ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0  ),
    ( 0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0  ),
    ( 0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0  ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0  ),
    ( 0,    -2,    -3,    -4,    -3,    -2,     0,     2,     3,     4,     3,     2,     0  ),
    ( 0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0  ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0  ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0  ),
    ( 0,    -2,    -3,    -4,    -3,    -2,     0,     2,     3,     4,     3,     2,     0  ),
    ( 0,     2,     3,     4,     3,     2,     0,    -2,    -3,    -4,    -3,    -2,     0  ),
    ( 0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0  ),
    ( 0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0  ),
    ( 0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0  ),
    ( 0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0  ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0  ),
    ( 0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0  ),
    ( 0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0  ),
    ( 0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0  ),
    ( 0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0  ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0  ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0  ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0  ),
    ( 0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0  ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0  ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0  ),
    ( 0,     2,     3,     4,     3,     2,     0,    -2,    -3,    -4,    -3,    -2,     0  ),
    ( 0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0  ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0  ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0  ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0  ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0  ),
    ( 0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0  ),
    ( 0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0  ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0  ),
    ( 0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0  ),
    ( 0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  )
    );

    Constant x2_sin_pairs : pairs_table := 
    -- x2 sin
    (
    ( 0,    -2,    -3,    -4,    -3,    -2,     0,     2,     3,     4,     3,     2,     0  ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0  ),
    ( 0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0  ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0  ),
    ( 0,    -2,    -3,    -4,    -3,    -2,     0,     2,     3,     4,     3,     2,     0  ),
    ( 0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0  ),
    ( 0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0  ),
    ( 0,     2,     3,     4,     3,     2,     0,    -2,    -3,    -4,    -3,    -2,     0  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0  ),
    ( 0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0  ),
    ( 0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0  ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0  ),
    ( 0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0  ),
    ( 0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0  ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0  ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0  ),
    ( 0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0  ),
    ( 0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0  ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0  ),
    ( 0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0  ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0  ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0  ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0  ),
    ( 0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0  ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0  ),
    ( 0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0  ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0  ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0  ),
    ( 0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0  ),
    ( 0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0  ),
    ( 0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0  ),
    ( 0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0  ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0  ),
    ( 0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0  ),
    ( 0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0  ),
    ( 0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0  ),
    ( 0,    -2,    -3,    -4,    -3,    -2,     0,     2,     3,     4,     3,     2,     0  ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0  ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0  ),
    ( 0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0  ),
    ( 0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0  ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0  ),
    ( 0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0  ),
    ( 0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0  )
    );

    Constant y2_cos_pairs : pairs_table := 
    -- y2 cos
    (
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3 ),
    ( 1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1  ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( 1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1  ),
    ( 1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1  ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2 ),
    ( 3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3  ),
    ( 3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3  ),
    ( 4,     3,     2,     0,    -2,    -3,    -4,    -3,    -2,     0,     2,     3,     4  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2 ),
    ( -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2 ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1  ),
    ( 3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3  ),
    ( 3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3  ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( -4,    -3,    -2,     0,     2,     3,     4,     3,     2,     0,    -2,    -3,    -4 ),
    ( -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2 ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( -4,    -3,    -2,     0,     2,     3,     4,     3,     2,     0,    -2,    -3,    -4 ),
    ( 4,     3,     2,     0,    -2,    -3,    -4,    -3,    -2,     0,     2,     3,     4  ),
    ( -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3 ),
    ( 3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3  ),
    ( 3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3  ),
    ( -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2 ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( 3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3  ),
    ( 3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3  ),
    ( 1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1  ),
    ( 1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1  ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( 3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3  ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( 4,     3,     2,     0,    -2,    -3,    -4,    -3,    -2,     0,     2,     3,     4  ),
    ( 3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3  ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( 3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3  ),
    ( 3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3  ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2 ),
    ( -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  )
    );
    
    Constant x2_cos_pairs : pairs_table := 
    -- x2 cos
    (
    ( -4,    -3,    -2,     0,     2,     3,     4,     3,     2,     0,    -2,    -3,    -4 ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( 1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1  ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( -4,    -3,    -2,     0,     2,     3,     4,     3,     2,     0,    -2,    -3,    -4 ),
    ( -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3 ),
    ( 1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1  ),
    ( 4,     3,     2,     0,    -2,    -3,    -4,    -3,    -2,     0,     2,     3,     4  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( 3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3  ),
    ( 1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1  ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2 ),
    ( 1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1  ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3 ),
    ( -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2 ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( 3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1  ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1  ),
    ( -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3 ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2 ),
    ( 1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1  ),
    ( -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3 ),
    ( -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3 ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3 ),
    ( -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3 ),
    ( 1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1  ),
    ( -4,    -3,    -2,     0,     2,     3,     4,     3,     2,     0,    -2,    -3,    -4 ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( 1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1  ),
    ( 3,     3,     2,     0,    -2,    -3,    -3,    -3,    -2,     0,     2,     3,     3  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( -2,    -2,    -1,     0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2 ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( 2,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,     2  ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( 1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1  ),
    ( 0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0  ),
    ( -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -1 ),
    ( -3,    -3,    -2,     0,     2,     3,     3,     3,     2,     0,    -2,    -3,    -3 )
    );
    

    --------------------------------------------------------- port map
    
    -- �⨤�� arctan(y/x)
    component cordic  
        port(
            clk : in STD_LOGIC;
            rst : in STD_LOGIC;
            x_in : in STD_LOGIC_VECTOR(14 downto 0);
            y_in : in STD_LOGIC_VECTOR(14 downto 0);
            x_out : out STD_LOGIC_VECTOR(17 downto 0);
            y_out : out STD_LOGIC_VECTOR(17 downto 0);
            z_out : out STD_LOGIC_VECTOR(7 downto 0)
        );
    end component;
    signal w_x_in : STD_LOGIC_VECTOR(14 downto 0);  ---
    signal w_y_in : STD_LOGIC_VECTOR(14 downto 0);
    COMPONENT ram_200x84
        PORT (
            clka : IN STD_LOGIC;
            wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
            addra : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
            dina : IN STD_LOGIC_VECTOR(83 DOWNTO 0);
            clkb : IN STD_LOGIC;
            addrb : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
            doutb : OUT STD_LOGIC_VECTOR(83 DOWNTO 0)
        );
    END COMPONENT;


    component ping_pong_buffer 
    port(
        clk : in std_logic;
        rst : in std_logic;	
        video_data:in std_logic_vector(7 downto 0);
        vga_hs_cnt :in integer range 0 to 857;	
        vga_vs_cnt :in integer range 0 to 524;
        ping_pong_out_8:out std_logic_vector(7 downto 0);
        ping_pong_out_7:out std_logic_vector(7 downto 0);
        ping_pong_out_6:out std_logic_vector(7 downto 0);
        ping_pong_out_5:out std_logic_vector(7 downto 0);
        ping_pong_out_4:out std_logic_vector(7 downto 0);
        ping_pong_out_3:out std_logic_vector(7 downto 0);
        ping_pong_out_2:out std_logic_vector(7 downto 0);
        ping_pong_out_1:out std_logic_vector(7 downto 0)
    );

    end component;


begin

ping_pong_out_2_out<=ping_pong_out_2;

--------------------------------------------------------- port map

  
ping_pong_buffer_0: ping_pong_buffer 
port map(
        clk 			=>clk 		     ,
        rst             =>rst            ,
		video_data      =>video_data     ,
		vga_hs_cnt      =>vga_hs_cnt     ,
		vga_vs_cnt      =>vga_vs_cnt     ,
		ping_pong_out_8 =>ping_pong_out_8,
		ping_pong_out_7 =>ping_pong_out_7,
		ping_pong_out_6 =>ping_pong_out_6,
		ping_pong_out_5 =>ping_pong_out_5,
		ping_pong_out_4 =>ping_pong_out_4,
		ping_pong_out_3 =>ping_pong_out_3,
		ping_pong_out_2 =>ping_pong_out_2,
		ping_pong_out_1 =>ping_pong_out_1
 );
 w_x_in <= std_logic_vector( abs(centroid_x_out) );
 w_y_in <= std_logic_vector( abs(centroid_y_out) );
cordic_1:cordic
port map(
		clk =>clk, 
		rst =>rst, 
		x_in => w_x_in,
		y_in => w_y_in, 
		x_out =>x_out,
		y_out =>y_out,	
		z_out =>z_out
);

--------------------------------------------------------- delay signal	
process(clk,rst)
begin
    if rst = '0' then
        kn_stage<=(others=>'0');
        
    elsif rising_edge(clk) then	
        kn_stage(0)<=kp_en;
        kn_stage(1)<=kn_stage(0);
        kn_stage(2)<=kn_stage(1);
        kn_stage(3)<=kn_stage(2);
        kn_stage(4)<=kn_stage(3);
        
        centroid_array_1<=centroid_array;
        centroid_array_2<=centroid_array_1;
        centroid_array_3<=centroid_array_2;
--        pepiclk<= 2 ;
    end if;
end process;

--------------------------------------------------------- line buffer
process(clk,rst)
begin
    if rst = '0' then
        centroid_array<=(others=>(others=>(others=>'0')));
    elsif rising_edge(clk) then
        centroid_array( 4, 4) <= ping_pong_out_8;
        centroid_array( 3, 4) <= ping_pong_out_7;
        centroid_array( 2, 4) <= ping_pong_out_6;
        centroid_array( 1, 4) <= ping_pong_out_5;
        centroid_array( 0, 4) <= ping_pong_out_4;
        centroid_array(-1, 4) <= ping_pong_out_3;
        centroid_array(-2, 4) <= ping_pong_out_2;
        centroid_array(-3, 4) <= ping_pong_out_1;
        centroid_array(-4, 4) <= video_data;
        
        centroid_array( 4, 3) <= centroid_array( 4, 4);
        centroid_array( 3, 3) <= centroid_array( 3, 4);
        centroid_array( 2, 3) <= centroid_array( 2, 4);
        centroid_array( 1, 3) <= centroid_array( 1, 4);
        centroid_array( 0, 3) <= centroid_array( 0, 4);
        centroid_array(-1, 3) <= centroid_array(-1, 4);
        centroid_array(-2, 3) <= centroid_array(-2, 4);
        centroid_array(-3, 3) <= centroid_array(-3, 4);
        centroid_array(-4, 3) <= centroid_array(-4, 4);
        
        centroid_array( 4, 2) <= centroid_array( 4, 3);
        centroid_array( 3, 2) <= centroid_array( 3, 3);
        centroid_array( 2, 2) <= centroid_array( 2, 3);
        centroid_array( 1, 2) <= centroid_array( 1, 3);
        centroid_array( 0, 2) <= centroid_array( 0, 3);
        centroid_array(-1, 2) <= centroid_array(-1, 3);
        centroid_array(-2, 2) <= centroid_array(-2, 3);
        centroid_array(-3, 2) <= centroid_array(-3, 3);
        centroid_array(-4, 2) <= centroid_array(-4, 3);
        
        centroid_array( 4, 1) <= centroid_array( 4, 2);
        centroid_array( 3, 1) <= centroid_array( 3, 2);
        centroid_array( 2, 1) <= centroid_array( 2, 2);
        centroid_array( 1, 1) <= centroid_array( 1, 2);
        centroid_array( 0, 1) <= centroid_array( 0, 2);
        centroid_array(-1, 1) <= centroid_array(-1, 2);
        centroid_array(-2, 1) <= centroid_array(-2, 2);
        centroid_array(-3, 1) <= centroid_array(-3, 2);
        centroid_array(-4, 1) <= centroid_array(-4, 2);
        
        centroid_array( 4, 0) <= centroid_array( 4, 1);
        centroid_array( 3, 0) <= centroid_array( 3, 1);
        centroid_array( 2, 0) <= centroid_array( 2, 1);
        centroid_array( 1, 0) <= centroid_array( 1, 1);
        centroid_array( 0, 0) <= centroid_array( 0, 1);
        centroid_array(-1, 0) <= centroid_array(-1, 1);
        centroid_array(-2, 0) <= centroid_array(-2, 1);
        centroid_array(-3, 0) <= centroid_array(-3, 1);
        centroid_array(-4, 0) <= centroid_array(-4, 1);
        
        centroid_array( 4,-1) <= centroid_array( 4, 0);
        centroid_array( 3,-1) <= centroid_array( 3, 0);
        centroid_array( 2,-1) <= centroid_array( 2, 0);
        centroid_array( 1,-1) <= centroid_array( 1, 0);
        centroid_array( 0,-1) <= centroid_array( 0, 0);
        centroid_array(-1,-1) <= centroid_array(-1, 0);
        centroid_array(-2,-1) <= centroid_array(-2, 0);
        centroid_array(-3,-1) <= centroid_array(-3, 0);
        centroid_array(-4,-1) <= centroid_array(-4, 0);
        
        centroid_array( 4,-2) <= centroid_array( 4,-1);
        centroid_array( 3,-2) <= centroid_array( 3,-1);
        centroid_array( 2,-2) <= centroid_array( 2,-1);
        centroid_array( 1,-2) <= centroid_array( 1,-1);
        centroid_array( 0,-2) <= centroid_array( 0,-1);
        centroid_array(-1,-2) <= centroid_array(-1,-1);
        centroid_array(-2,-2) <= centroid_array(-2,-1);
        centroid_array(-3,-2) <= centroid_array(-3,-1);
        centroid_array(-4,-2) <= centroid_array(-4,-1);
        
        centroid_array( 4,-3) <= centroid_array( 4,-2);
        centroid_array( 3,-3) <= centroid_array( 3,-2);
        centroid_array( 2,-3) <= centroid_array( 2,-2);
        centroid_array( 1,-3) <= centroid_array( 1,-2);
        centroid_array( 0,-3) <= centroid_array( 0,-2);
        centroid_array(-1,-3) <= centroid_array(-1,-2);
        centroid_array(-2,-3) <= centroid_array(-2,-2);
        centroid_array(-3,-3) <= centroid_array(-3,-2);
        centroid_array(-4,-3) <= centroid_array(-4,-2);
        
        centroid_array( 4,-4) <= centroid_array( 4,-3);
        centroid_array( 3,-4) <= centroid_array( 3,-3);
        centroid_array( 2,-4) <= centroid_array( 2,-3);
        centroid_array( 1,-4) <= centroid_array( 1,-3);
        centroid_array( 0,-4) <= centroid_array( 0,-3);
        centroid_array(-1,-4) <= centroid_array(-1,-3);
        centroid_array(-2,-4) <= centroid_array(-2,-3);
        centroid_array(-3,-4) <= centroid_array(-3,-3);
        centroid_array(-4,-4) <= centroid_array(-4,-3);
--        pepiclk<= 3 ;
    end if;
end process;

--------------------------------------------------------- Sobel �j�׭p��
process(clk,rst)
    variable centroid_x:signed(14 downto 0):=(others=>'0');
    variable centroid_y:signed(14 downto 0):=(others=>'0');
begin

if rst = '0' then
	centroid_x_out <= (others=>'0');
	centroid_y_out <= (others=>'0');
--	pepiclk<= 4 ;
elsif rising_edge(clk) then
	centroid_x:=(others=>'0');
	centroid_y:=(others=>'0');
    
--centroid_array is from ORB_result
	for step in -4 to 4 loop
        centroid_x := centroid_x - resize(signed('0'  &centroid_array(step,-4)&'0'),15 ) 
                                 - resize(signed("00" &centroid_array(step,-3)+centroid_array(step,-3)(7 downto 1)),15 )
                                 - resize(signed('0'  &centroid_array(step,-2)),15 )
                                 - resize(signed('0'  &centroid_array(step,-1)(7 downto 1)),15 )
                                 + resize(signed('0'  &centroid_array(step,1)(7 downto 1)),15 )
                                 + resize(signed('0'  &centroid_array(step,2)),15 )
                                 + resize(signed("00" &centroid_array(step,3)+centroid_array(step,3)(7 downto 1)),15 )
                                 + resize(signed('0'  &centroid_array(step,4)&'0'),15 );
                                                      
        centroid_y := centroid_y - resize(signed('0'  &centroid_array(-4,step)&'0'),15 )
                                 - resize(signed("00" &centroid_array(-3,step) + centroid_array(-3,step)(7 downto 1)),15 )
                                 - resize(signed('0'  &centroid_array(-2,step)),15 )
                                 - resize(signed('0'  &centroid_array(-1,step)(7 downto 1)),15 )
                                 + resize(signed('0'  &centroid_array(1,step)(7 downto 1)),15 )
                                 + resize(signed('0'  &centroid_array(2,step)),15 )
                                 + resize(signed("00" &centroid_array(3,step) + centroid_array(3,step)(7 downto 1)),15 )
                                 + resize(signed('0'  &centroid_array(4,step)&'0'),15 );
	end loop;
    
	centroid_y_out <= centroid_y;	
	centroid_x_out <= centroid_x; 
	
end if;
end process;

--------------------------------------------------------- ���׭p��

process(rst, clk )
begin
    if rst='0' then
        centroid_angle <= 0 ;
    elsif rising_edge(clk)then
        
        if    (centroid_x_out(14) = '0' and centroid_y_out(14) = '0')then --��1�H��  
            centroid_angle <= 000 + conv_integer(z_out);
            --            pepiclk<= 5 ;
        elsif (centroid_x_out(14) = '1' and centroid_y_out(14) = '0')then --��2�H��  
            centroid_angle <= 180 - conv_integer(z_out);
            
        elsif (centroid_x_out(14) = '1' and centroid_y_out(14) = '1')then --��3�H��  
            centroid_angle <= 180 + conv_integer(z_out);
            
        elsif (centroid_x_out(14) = '0' and centroid_y_out(14) = '1')then --��4�H��  
            centroid_angle <= 360 - conv_integer(z_out);
            
        end if;
        
    end if;
end process;

--after centroid_array has been process with cordic
process(rst, clk )
begin
    if rst='0'then
        angle_range<=0;	
    elsif rising_edge(clk)then
	
           if (centroid_angle< 15	or  centroid_angle >= 345) then		angle_range <= 0;
        elsif (centroid_angle< 45	and centroid_angle >= 15 ) then		angle_range <= 1;
        elsif (centroid_angle< 75	and centroid_angle >= 45 ) then		angle_range <= 2;
        elsif (centroid_angle< 105	and centroid_angle >= 75 ) then		angle_range <= 3;
        elsif (centroid_angle< 135	and centroid_angle >= 105) then		angle_range <= 4;
        elsif (centroid_angle< 165	and centroid_angle >= 135) then		angle_range <= 5;
        elsif (centroid_angle< 195	and centroid_angle >= 165) then		angle_range <= 6;
        elsif (centroid_angle< 225	and centroid_angle >= 195) then		angle_range <= 7;
        elsif (centroid_angle< 255	and centroid_angle >= 225) then		angle_range <= 8;
        elsif (centroid_angle< 285	and centroid_angle >= 255) then		angle_range <= 9;
        elsif (centroid_angle< 315	and centroid_angle >= 285) then		angle_range <= 10;
        elsif (centroid_angle< 345	and centroid_angle >= 315) then		angle_range <= 11;
--        pepiclk<= 6 ;
        end if;

    end if;
end process;

--------------------------------------------------------- brief calculate
process(clk,rst)
    variable steered_y_1    :integer range -9 to 9;
    variable steered_x_1    :integer range -9 to 9;
    variable steered_y_2    :integer range -9 to 9;
    variable steered_x_2    :integer range -9 to 9;
    
    variable steered_y_1_for_kerenl    :integer range -4 to 4;
    variable steered_x_1_for_kerenl    :integer range -4 to 4;
    variable steered_y_2_for_kerenl    :integer range -4 to 4;
    variable steered_x_2_for_kerenl    :integer range -4 to 4;
    
begin
    if rst='0'then
        brief_code<=(others=>'0');
    elsif rising_edge(clk)then

        for pair in 0 to (pairs_num-1) loop --    pairs_num : integer:=64;
            -- y' = sin(�c) * x + cos(�c) * y
            -- x' = cos(�c) * x - sin(�c) * y
            
            steered_y_1 := x1_sin_pairs(pair, angle_range) + y1_cos_pairs(pair, angle_range);
            steered_x_1 := x1_cos_pairs(pair, angle_range) - y1_sin_pairs(pair, angle_range);
            
            steered_y_2 := x2_sin_pairs(pair, angle_range) + y2_cos_pairs(pair, angle_range);
            steered_x_2 := x2_cos_pairs(pair, angle_range) - y2_sin_pairs(pair, angle_range);
            
            if -5 > steered_y_1 then
                steered_y_1_for_kerenl := -4;
            elsif steered_y_1 > 5  then
                steered_y_1_for_kerenl :=  4;
            else 
                steered_y_1_for_kerenl := steered_y_1;
            end if ;
            
            if -5 > steered_x_1 then
                steered_x_1_for_kerenl := -4;
            elsif steered_x_1 > 5  then
                steered_x_1_for_kerenl :=  4;
            else 
                steered_x_1_for_kerenl := steered_x_1;
            end if ;
            
            if -5 > steered_y_2 then
                steered_y_2_for_kerenl := -4;
            elsif steered_y_2 > 5  then
                steered_y_2_for_kerenl :=  4;
            else 
                steered_y_2_for_kerenl := steered_y_2;
            end if ;
            
            if -5 > steered_x_2 then
                steered_x_2_for_kerenl := -4;
            elsif steered_x_2 > 5  then
                steered_x_2_for_kerenl :=  4;
            else 
                steered_x_2_for_kerenl := steered_x_2;
            end if ;
            
            
            if centroid_array_3( steered_y_1_for_kerenl , steered_x_1_for_kerenl ) > centroid_array_3( steered_y_2_for_kerenl , steered_x_2_for_kerenl )then
                brief_code(pair) <='1';
--                pepiclk<= 8 ;
            else
                brief_code(pair) <='0';
            end if;
            
        end loop;


    end if;
end process;

--------------------------------------------------------------------------------------
--------------------------------------------------------- save data
process(clk,rst)
begin
if rst='0'then

BOUT_1  <= (others=>'0');
elsif rising_edge(clk)then

----------------trak---------
--        if rising_edge(video_clk) then
--            if (vga_hs_cnt > TRACKX - TRACKSQ  and vga_hs_cnt < TRACKX + TRACKSQ
--	        and vga_vs_cnt > TRACKY - TRACKSQ  and vga_vs_cnt < TRACKY + TRACKSQ
--	     	and vga_hs_cnt > 64 and vga_hs_cnt < 656
--	        and vga_vs_cnt > 32 and vga_vs_cnt < 448      ) then
---------------------------------------------------------    
		--image 1
		if (vga_hs_cnt > 0  and vga_hs_cnt < 720 
	and vga_vs_cnt>= 0 and vga_vs_cnt< 480 ) then
			if kn_stage(4)='1' then
                BOUT_1  <= brief_code & std_logic_vector(to_unsigned(vga_vs_cnt,10)) & std_logic_vector(to_unsigned(vga_hs_cnt,10));
--                pepiclk<= 9 ;
		end if;
       end if;

end if;
end process;
end Behavioral;	